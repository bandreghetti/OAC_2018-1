library verilog;
use verilog.vl_types.all;
entity Subtrator_vlg_vec_tst is
end Subtrator_vlg_vec_tst;
