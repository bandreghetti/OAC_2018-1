Mux8_inst : Mux8 PORT MAP (
		data0	 => data0_sig,
		data1	 => data1_sig,
		data2	 => data2_sig,
		data3	 => data3_sig,
		data4	 => data4_sig,
		data5	 => data5_sig,
		data6	 => data6_sig,
		data7	 => data7_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
