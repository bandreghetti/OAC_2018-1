library verilog;
use verilog.vl_types.all;
entity Controlador_vlg_vec_tst is
end Controlador_vlg_vec_tst;
