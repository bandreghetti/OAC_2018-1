library verilog;
use verilog.vl_types.all;
entity Somador_vlg_check_tst is
    port(
        C_out           : in     vl_logic;
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Somador_vlg_check_tst;
