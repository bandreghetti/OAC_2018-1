library verilog;
use verilog.vl_types.all;
entity RegBank_vlg_vec_tst is
end RegBank_vlg_vec_tst;
