Mux4_inst : Mux4 PORT MAP (
		data0	 => data0_sig,
		data1	 => data1_sig,
		data2	 => data2_sig,
		data3	 => data3_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
