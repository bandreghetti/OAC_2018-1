library verilog;
use verilog.vl_types.all;
entity ULA_32bits_vlg_vec_tst is
end ULA_32bits_vlg_vec_tst;
