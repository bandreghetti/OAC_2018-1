library verilog;
use verilog.vl_types.all;
entity reg32_vlg_vec_tst is
end reg32_vlg_vec_tst;
