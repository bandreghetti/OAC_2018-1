library verilog;
use verilog.vl_types.all;
entity Somador_vlg_vec_tst is
end Somador_vlg_vec_tst;
