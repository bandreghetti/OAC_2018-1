library verilog;
use verilog.vl_types.all;
entity ULA_Full_vlg_vec_tst is
end ULA_Full_vlg_vec_tst;
